LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity BIT4fulladder is
    Port ( A0,A1,A2,A3,B0,B1,B2,B3 : in  STD_LOGIC;
           CIN : in  STD_LOGIC;
           S0,S1,S2,S3 : out  STD_LOGIC;
           CARRY : out  STD_LOGIC);
end BIT4fulladder;
architecture Behavioral of BIT4fulladder is
SIGNAL C1,C2,C3:STD_LOGIC;
COMPONENT BITFULLADDER
PORT(A,B,CIN:IN STD_LOGIC;SUM,CARRY:OUT STD_LOGIC);
END COMPONENT;
begin
STEP7:BITFULLADDER PORT MAP(A0,B0,CIN,S0,C1);
STEP8:BITFULLADDER PORT MAP(A1,B1,C1,S1,C2);
STEP9:BITFULLADDER PORT MAP(A2,B2,C2,S2,C3);
STEP10:BITFULLADDER PORT MAP(A3,B3,C3,S3,CARRY);
end Behavioral;